 module tb;

    // Inputs
    reg [6271:0] A;
    reg [71:0] B;
    // Outputs
    wire [5407:0] Res;

    // Instantiate the Unit Under Test (UUT)
    e_Mat_mult uut (
        .A(A), 
        .B(B), 
        .Res(Res)
    );

    initial begin
        // Apply Inputs
        A = 0;  B = 0;  #100;
        B = {8'd1,8'd2,8'd3,8'd4,8'd5,8'd6,8'd7,8'd8,8'd9};
        A = {8'd10,8'd11,8'd12,8'd13,8'd14,8'd15,8'd16,8'd17,8'd18,8'd19,8'd20,8'd21,8'd22,8'd23,8'd24,8'd25,8'd26,8'd27,8'd28,8'd29,8'd30,8'd31,8'd32,8'd33,8'd34,8'd35,8'd36,8'd37,8'd38,8'd39,8'd40,8'd41,8'd42,8'd43,8'd44,8'd45,8'd46,8'd47,8'd48,8'd49,8'd50,8'd51,8'd52,8'd53,8'd54,8'd55,8'd56,8'd57,8'd58,8'd59,8'd60,8'd61,8'd62,8'd63,8'd64,8'd65,8'd66,8'd67,8'd68,8'd69,8'd70,8'd71,8'd72,8'd73,8'd74,8'd75,8'd76,8'd77,8'd78,8'd79,8'd80,8'd81,8'd82,8'd83,8'd84,8'd85,8'd86,8'd87,8'd88,8'd89,8'd90,8'd91,8'd92,8'd93,8'd94,8'd95,8'd96,8'd97,8'd98,8'd99,8'd100,8'd101,8'd102,8'd103,8'd104,8'd105,8'd106,8'd107,8'd108,8'd109,8'd110,8'd111,8'd112,8'd113,8'd114,8'd115,8'd116,8'd117,8'd118,8'd119,8'd120,8'd121,8'd122,8'd123,8'd124,8'd125,8'd126,8'd127,8'd128,8'd129,8'd130,8'd131,8'd132,8'd133,8'd134,8'd135,8'd136,8'd137,8'd138,8'd139,8'd140,8'd141,8'd142,8'd143,8'd144,8'd145,8'd146,8'd147,8'd148,8'd149,8'd150,8'd151,8'd152,8'd153,8'd154,8'd155,8'd156,8'd157,8'd158,8'd159,8'd160,8'd161,8'd162,8'd163,8'd164,8'd165,8'd166,8'd167,8'd168,8'd169,8'd170,8'd171,8'd172,8'd173,8'd174,8'd175,8'd176,8'd177,8'd178,8'd179,8'd180,8'd181,8'd182,8'd183,8'd184,8'd185,8'd186,8'd187,8'd188,8'd189,8'd190,8'd191,8'd192,8'd193,8'd194,8'd195,8'd196,8'd197,8'd198,8'd199,8'd200,8'd201,8'd202,8'd203,8'd204,8'd205,8'd206,8'd207,8'd208,8'd209,8'd210,8'd211,8'd212,8'd213,8'd214,8'd215,8'd216,8'd217,8'd218,8'd219,8'd220,8'd221,8'd222,8'd223,8'd224,8'd225,8'd226,8'd227,8'd228,8'd229,8'd230,8'd231,8'd232,8'd233,8'd234,8'd235,8'd236,8'd237,8'd238,8'd239,8'd240,8'd241,8'd242,8'd243,8'd244,8'd245,8'd246,8'd247,8'd248,8'd249,8'd250,8'd251,8'd252,8'd253,8'd254,8'd255,8'd256,8'd257,8'd258,8'd259,8'd260,8'd261,8'd262,8'd263,8'd264,8'd265,8'd266,8'd267,8'd268,8'd269,8'd270,8'd271,8'd272,8'd273,8'd274,8'd275,8'd276,8'd277,8'd278,8'd279,8'd280,8'd281,8'd282,8'd283,8'd284,8'd285,8'd286,8'd287,8'd288,8'd289,8'd290,8'd291,8'd292,8'd293,8'd294,8'd295,8'd296,8'd297,8'd298,8'd299,8'd300,8'd301,8'd302,8'd303,8'd304,8'd305,8'd306,8'd307,8'd308,8'd309,8'd310,8'd311,8'd312,8'd313,8'd314,8'd315,8'd316,8'd317,8'd318,8'd319,8'd320,8'd321,8'd322,8'd323,8'd324,8'd325,8'd326,8'd327,8'd328,8'd329,8'd330,8'd331,8'd332,8'd333,8'd334,8'd335,8'd336,8'd337,8'd338,8'd339,8'd340,8'd341,8'd342,8'd343,8'd344,8'd345,8'd346,8'd347,8'd348,8'd349,8'd350,8'd351,8'd352,8'd353,8'd354,8'd355,8'd356,8'd357,8'd358,8'd359,8'd360,8'd361,8'd362,8'd363,8'd364,8'd365,8'd366,8'd367,8'd368,8'd369,8'd370,8'd371,8'd372,8'd373,8'd374,8'd375,8'd376,8'd377,8'd378,8'd379,8'd380,8'd381,8'd382,8'd383,8'd384,8'd385,8'd386,8'd387,8'd388,8'd389,8'd390,8'd391,8'd392,8'd393,8'd394,8'd395,8'd396,8'd397,8'd398,8'd399,8'd400,8'd401,8'd402,8'd403,8'd404,8'd405,8'd406,8'd407,8'd408,8'd409,8'd410,8'd411,8'd412,8'd413,8'd414,8'd415,8'd416,8'd417,8'd418,8'd419,8'd420,8'd421,8'd422,8'd423,8'd424,8'd425,8'd426,8'd427,8'd428,8'd429,8'd430,8'd431,8'd432,8'd433,8'd434,8'd435,8'd436,8'd437,8'd438,8'd439,8'd440,8'd441,8'd442,8'd443,8'd444,8'd445,8'd446,8'd447,8'd448,8'd449,8'd450,8'd451,8'd452,8'd453,8'd454,8'd455,8'd456,8'd457,8'd458,8'd459,8'd460,8'd461,8'd462,8'd463,8'd464,8'd465,8'd466,8'd467,8'd468,8'd469,8'd470,8'd471,8'd472,8'd473,8'd474,8'd475,8'd476,8'd477,8'd478,8'd479,8'd480,8'd481,8'd482,8'd483,8'd484,8'd485,8'd486,8'd487,8'd488,8'd489,8'd490,8'd491,8'd492,8'd493,8'd494,8'd495,8'd496,8'd497,8'd498,8'd499,8'd500,8'd501,8'd502,8'd503,8'd504,8'd505,8'd506,8'd507,8'd508,8'd509,8'd510,8'd511,8'd512,8'd513,8'd514,8'd515,8'd516,8'd517,8'd518,8'd519,8'd520,8'd521,8'd522,8'd523,8'd524,8'd525,8'd526,8'd527,8'd528,8'd529,8'd530,8'd531,8'd532,8'd533,8'd534,8'd535,8'd536,8'd537,8'd538,8'd539,8'd540,8'd541,8'd542,8'd543,8'd544,8'd545,8'd546,8'd547,8'd548,8'd549,8'd550,8'd551,8'd552,8'd553,8'd554,8'd555,8'd556,8'd557,8'd558,8'd559,8'd560,8'd561,8'd562,8'd563,8'd564,8'd565,8'd566,8'd567,8'd568,8'd569,8'd570,8'd571,8'd572,8'd573,8'd574,8'd575,8'd576,8'd577,8'd578,8'd579,8'd580,8'd581,8'd582,8'd583,8'd584,8'd585,8'd586,8'd587,8'd588,8'd589,8'd590,8'd591,8'd592,8'd593,8'd594,8'd595,8'd596,8'd597,8'd598,8'd599,8'd600,8'd601,8'd602,8'd603,8'd604,8'd605,8'd606,8'd607,8'd608,8'd609,8'd610,8'd611,8'd612,8'd613,8'd614,8'd615,8'd616,8'd617,8'd618,8'd619,8'd620,8'd621,8'd622,8'd623,8'd624,8'd625,8'd626,8'd627,8'd628,8'd629,8'd630,8'd631,8'd632,8'd633,8'd634,8'd635,8'd636,8'd637,8'd638,8'd639,8'd640,8'd641,8'd642,8'd643,8'd644,8'd645,8'd646,8'd647,8'd648,8'd649,8'd650,8'd651,8'd652,8'd653,8'd654,8'd655,8'd656,8'd657,8'd658,8'd659,8'd660,8'd661,8'd662,8'd663,8'd664,8'd665,8'd666,8'd667,8'd668,8'd669,8'd670,8'd671,8'd672,8'd673,8'd674,8'd675,8'd676,8'd677,8'd678,8'd679,8'd680,8'd681,8'd682,8'd683,8'd684,8'd685,8'd686,8'd687,8'd688,8'd689,8'd690,8'd691,8'd692,8'd693,8'd694,8'd695,8'd696,8'd697,8'd698,8'd699,8'd700,8'd701,8'd702,8'd703,8'd704,8'd705,8'd706,8'd707,8'd708,8'd709,8'd710,8'd711,8'd712,8'd713,8'd714,8'd715,8'd716,8'd717,8'd718,8'd719,8'd720,8'd721,8'd722,8'd723,8'd724,8'd725,8'd726,8'd727,8'd728,8'd729,8'd730,8'd731,8'd732,8'd733,8'd734,8'd735,8'd736,8'd737,8'd738,8'd739,8'd740,8'd741,8'd742,8'd743,8'd744,8'd745,8'd746,8'd747,8'd748,8'd749,8'd750,8'd751,8'd752,8'd753,8'd754,8'd755,8'd756,8'd757,8'd758,8'd759,8'd760,8'd761,8'd762,8'd763,8'd764,8'd765,8'd766,8'd767,8'd768,8'd769,8'd770,8'd771,8'd772,8'd773,8'd774,8'd775,8'd776,8'd777,8'd778,8'd779,8'd780,8'd781,8'd782,8'd783,8'd784,8'd785,8'd786,8'd787,8'd788,8'd789,8'd790,8'd791,8'd792,8'd793};
    end
      
endmodule