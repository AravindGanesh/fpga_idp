 //Module for applying Sobel filter on a 28x28 image
//Where A is 28x28 matrix and B is 3x3 matrix
module sobel_filter(A,B,Res);
    
    //input and output ports.
    //input clk;
    //The size 6272 bits which is 28*28=784 elements,each of which is 5 bits wide.    
    input [3919:0] A;
    //The size 27 bits which is 3*3=9 elements,each of which is 3 bits wide.
    input [26:0] B;
    //The size 5408 bits which is 26*26=676 elements,each of which is 8 bits wide.
    output [5407:0] Res;
    //internal variables 
    reg [5407:0] Res;
    reg [4:0] A1 [0:27][0:27];
    reg [2:0] B1 [0:2][0:2];
    reg [7:0] Res1 [0:25][0:25]; 
    integer i,j,k;

    //always @(negedge clk) begin
    initial begin
    //Initialize the matrices-convert 1 D to 3D arrays
        {A1[0][0],A1[0][1],A1[0][2],A1[0][3],A1[0][4],A1[0][5],A1[0][6],A1[0][7],A1[0][8],A1[0][9],A1[0][10],A1[0][11],A1[0][12],A1[0][13],A1[0][14],A1[0][15],A1[0][16],A1[0][17],A1[0][18],A1[0][19],A1[0][20],A1[0][21],A1[0][22],A1[0][23],A1[0][24],A1[0][25],A1[0][26],A1[0][27],A1[1][0],A1[1][1],A1[1][2],A1[1][3],A1[1][4],A1[1][5],A1[1][6],A1[1][7],A1[1][8],A1[1][9],A1[1][10],A1[1][11],A1[1][12],A1[1][13],A1[1][14],A1[1][15],A1[1][16],A1[1][17],A1[1][18],A1[1][19],A1[1][20],A1[1][21],A1[1][22],A1[1][23],A1[1][24],A1[1][25],A1[1][26],A1[1][27],A1[2][0],A1[2][1],A1[2][2],A1[2][3],A1[2][4],A1[2][5],A1[2][6],A1[2][7],A1[2][8],A1[2][9],A1[2][10],A1[2][11],A1[2][12],A1[2][13],A1[2][14],A1[2][15],A1[2][16],A1[2][17],A1[2][18],A1[2][19],A1[2][20],A1[2][21],A1[2][22],A1[2][23],A1[2][24],A1[2][25],A1[2][26],A1[2][27],A1[3][0],A1[3][1],A1[3][2],A1[3][3],A1[3][4],A1[3][5],A1[3][6],A1[3][7],A1[3][8],A1[3][9],A1[3][10],A1[3][11],A1[3][12],A1[3][13],A1[3][14],A1[3][15],A1[3][16],A1[3][17],A1[3][18],A1[3][19],A1[3][20],A1[3][21],A1[3][22],A1[3][23],A1[3][24],A1[3][25],A1[3][26],A1[3][27],A1[4][0],A1[4][1],A1[4][2],A1[4][3],A1[4][4],A1[4][5],A1[4][6],A1[4][7],A1[4][8],A1[4][9],A1[4][10],A1[4][11],A1[4][12],A1[4][13],A1[4][14],A1[4][15],A1[4][16],A1[4][17],A1[4][18],A1[4][19],A1[4][20],A1[4][21],A1[4][22],A1[4][23],A1[4][24],A1[4][25],A1[4][26],A1[4][27],A1[5][0],A1[5][1],A1[5][2],A1[5][3],A1[5][4],A1[5][5],A1[5][6],A1[5][7],A1[5][8],A1[5][9],A1[5][10],A1[5][11],A1[5][12],A1[5][13],A1[5][14],A1[5][15],A1[5][16],A1[5][17],A1[5][18],A1[5][19],A1[5][20],A1[5][21],A1[5][22],A1[5][23],A1[5][24],A1[5][25],A1[5][26],A1[5][27],A1[6][0],A1[6][1],A1[6][2],A1[6][3],A1[6][4],A1[6][5],A1[6][6],A1[6][7],A1[6][8],A1[6][9],A1[6][10],A1[6][11],A1[6][12],A1[6][13],A1[6][14],A1[6][15],A1[6][16],A1[6][17],A1[6][18],A1[6][19],A1[6][20],A1[6][21],A1[6][22],A1[6][23],A1[6][24],A1[6][25],A1[6][26],A1[6][27],A1[7][0],A1[7][1],A1[7][2],A1[7][3],A1[7][4],A1[7][5],A1[7][6],A1[7][7],A1[7][8],A1[7][9],A1[7][10],A1[7][11],A1[7][12],A1[7][13],A1[7][14],A1[7][15],A1[7][16],A1[7][17],A1[7][18],A1[7][19],A1[7][20],A1[7][21],A1[7][22],A1[7][23],A1[7][24],A1[7][25],A1[7][26],A1[7][27],A1[8][0],A1[8][1],A1[8][2],A1[8][3],A1[8][4],A1[8][5],A1[8][6],A1[8][7],A1[8][8],A1[8][9],A1[8][10],A1[8][11],A1[8][12],A1[8][13],A1[8][14],A1[8][15],A1[8][16],A1[8][17],A1[8][18],A1[8][19],A1[8][20],A1[8][21],A1[8][22],A1[8][23],A1[8][24],A1[8][25],A1[8][26],A1[8][27],A1[9][0],A1[9][1],A1[9][2],A1[9][3],A1[9][4],A1[9][5],A1[9][6],A1[9][7],A1[9][8],A1[9][9],A1[9][10],A1[9][11],A1[9][12],A1[9][13],A1[9][14],A1[9][15],A1[9][16],A1[9][17],A1[9][18],A1[9][19],A1[9][20],A1[9][21],A1[9][22],A1[9][23],A1[9][24],A1[9][25],A1[9][26],A1[9][27],A1[10][0],A1[10][1],A1[10][2],A1[10][3],A1[10][4],A1[10][5],A1[10][6],A1[10][7],A1[10][8],A1[10][9],A1[10][10],A1[10][11],A1[10][12],A1[10][13],A1[10][14],A1[10][15],A1[10][16],A1[10][17],A1[10][18],A1[10][19],A1[10][20],A1[10][21],A1[10][22],A1[10][23],A1[10][24],A1[10][25],A1[10][26],A1[10][27],A1[11][0],A1[11][1],A1[11][2],A1[11][3],A1[11][4],A1[11][5],A1[11][6],A1[11][7],A1[11][8],A1[11][9],A1[11][10],A1[11][11],A1[11][12],A1[11][13],A1[11][14],A1[11][15],A1[11][16],A1[11][17],A1[11][18],A1[11][19],A1[11][20],A1[11][21],A1[11][22],A1[11][23],A1[11][24],A1[11][25],A1[11][26],A1[11][27],A1[12][0],A1[12][1],A1[12][2],A1[12][3],A1[12][4],A1[12][5],A1[12][6],A1[12][7],A1[12][8],A1[12][9],A1[12][10],A1[12][11],A1[12][12],A1[12][13],A1[12][14],A1[12][15],A1[12][16],A1[12][17],A1[12][18],A1[12][19],A1[12][20],A1[12][21],A1[12][22],A1[12][23],A1[12][24],A1[12][25],A1[12][26],A1[12][27],A1[13][0],A1[13][1],A1[13][2],A1[13][3],A1[13][4],A1[13][5],A1[13][6],A1[13][7],A1[13][8],A1[13][9],A1[13][10],A1[13][11],A1[13][12],A1[13][13],A1[13][14],A1[13][15],A1[13][16],A1[13][17],A1[13][18],A1[13][19],A1[13][20],A1[13][21],A1[13][22],A1[13][23],A1[13][24],A1[13][25],A1[13][26],A1[13][27],A1[14][0],A1[14][1],A1[14][2],A1[14][3],A1[14][4],A1[14][5],A1[14][6],A1[14][7],A1[14][8],A1[14][9],A1[14][10],A1[14][11],A1[14][12],A1[14][13],A1[14][14],A1[14][15],A1[14][16],A1[14][17],A1[14][18],A1[14][19],A1[14][20],A1[14][21],A1[14][22],A1[14][23],A1[14][24],A1[14][25],A1[14][26],A1[14][27],A1[15][0],A1[15][1],A1[15][2],A1[15][3],A1[15][4],A1[15][5],A1[15][6],A1[15][7],A1[15][8],A1[15][9],A1[15][10],A1[15][11],A1[15][12],A1[15][13],A1[15][14],A1[15][15],A1[15][16],A1[15][17],A1[15][18],A1[15][19],A1[15][20],A1[15][21],A1[15][22],A1[15][23],A1[15][24],A1[15][25],A1[15][26],A1[15][27],A1[16][0],A1[16][1],A1[16][2],A1[16][3],A1[16][4],A1[16][5],A1[16][6],A1[16][7],A1[16][8],A1[16][9],A1[16][10],A1[16][11],A1[16][12],A1[16][13],A1[16][14],A1[16][15],A1[16][16],A1[16][17],A1[16][18],A1[16][19],A1[16][20],A1[16][21],A1[16][22],A1[16][23],A1[16][24],A1[16][25],A1[16][26],A1[16][27],A1[17][0],A1[17][1],A1[17][2],A1[17][3],A1[17][4],A1[17][5],A1[17][6],A1[17][7],A1[17][8],A1[17][9],A1[17][10],A1[17][11],A1[17][12],A1[17][13],A1[17][14],A1[17][15],A1[17][16],A1[17][17],A1[17][18],A1[17][19],A1[17][20],A1[17][21],A1[17][22],A1[17][23],A1[17][24],A1[17][25],A1[17][26],A1[17][27],A1[18][0],A1[18][1],A1[18][2],A1[18][3],A1[18][4],A1[18][5],A1[18][6],A1[18][7],A1[18][8],A1[18][9],A1[18][10],A1[18][11],A1[18][12],A1[18][13],A1[18][14],A1[18][15],A1[18][16],A1[18][17],A1[18][18],A1[18][19],A1[18][20],A1[18][21],A1[18][22],A1[18][23],A1[18][24],A1[18][25],A1[18][26],A1[18][27],A1[19][0],A1[19][1],A1[19][2],A1[19][3],A1[19][4],A1[19][5],A1[19][6],A1[19][7],A1[19][8],A1[19][9],A1[19][10],A1[19][11],A1[19][12],A1[19][13],A1[19][14],A1[19][15],A1[19][16],A1[19][17],A1[19][18],A1[19][19],A1[19][20],A1[19][21],A1[19][22],A1[19][23],A1[19][24],A1[19][25],A1[19][26],A1[19][27],A1[20][0],A1[20][1],A1[20][2],A1[20][3],A1[20][4],A1[20][5],A1[20][6],A1[20][7],A1[20][8],A1[20][9],A1[20][10],A1[20][11],A1[20][12],A1[20][13],A1[20][14],A1[20][15],A1[20][16],A1[20][17],A1[20][18],A1[20][19],A1[20][20],A1[20][21],A1[20][22],A1[20][23],A1[20][24],A1[20][25],A1[20][26],A1[20][27],A1[21][0],A1[21][1],A1[21][2],A1[21][3],A1[21][4],A1[21][5],A1[21][6],A1[21][7],A1[21][8],A1[21][9],A1[21][10],A1[21][11],A1[21][12],A1[21][13],A1[21][14],A1[21][15],A1[21][16],A1[21][17],A1[21][18],A1[21][19],A1[21][20],A1[21][21],A1[21][22],A1[21][23],A1[21][24],A1[21][25],A1[21][26],A1[21][27],A1[22][0],A1[22][1],A1[22][2],A1[22][3],A1[22][4],A1[22][5],A1[22][6],A1[22][7],A1[22][8],A1[22][9],A1[22][10],A1[22][11],A1[22][12],A1[22][13],A1[22][14],A1[22][15],A1[22][16],A1[22][17],A1[22][18],A1[22][19],A1[22][20],A1[22][21],A1[22][22],A1[22][23],A1[22][24],A1[22][25],A1[22][26],A1[22][27],A1[23][0],A1[23][1],A1[23][2],A1[23][3],A1[23][4],A1[23][5],A1[23][6],A1[23][7],A1[23][8],A1[23][9],A1[23][10],A1[23][11],A1[23][12],A1[23][13],A1[23][14],A1[23][15],A1[23][16],A1[23][17],A1[23][18],A1[23][19],A1[23][20],A1[23][21],A1[23][22],A1[23][23],A1[23][24],A1[23][25],A1[23][26],A1[23][27],A1[24][0],A1[24][1],A1[24][2],A1[24][3],A1[24][4],A1[24][5],A1[24][6],A1[24][7],A1[24][8],A1[24][9],A1[24][10],A1[24][11],A1[24][12],A1[24][13],A1[24][14],A1[24][15],A1[24][16],A1[24][17],A1[24][18],A1[24][19],A1[24][20],A1[24][21],A1[24][22],A1[24][23],A1[24][24],A1[24][25],A1[24][26],A1[24][27],A1[25][0],A1[25][1],A1[25][2],A1[25][3],A1[25][4],A1[25][5],A1[25][6],A1[25][7],A1[25][8],A1[25][9],A1[25][10],A1[25][11],A1[25][12],A1[25][13],A1[25][14],A1[25][15],A1[25][16],A1[25][17],A1[25][18],A1[25][19],A1[25][20],A1[25][21],A1[25][22],A1[25][23],A1[25][24],A1[25][25],A1[25][26],A1[25][27],A1[26][0],A1[26][1],A1[26][2],A1[26][3],A1[26][4],A1[26][5],A1[26][6],A1[26][7],A1[26][8],A1[26][9],A1[26][10],A1[26][11],A1[26][12],A1[26][13],A1[26][14],A1[26][15],A1[26][16],A1[26][17],A1[26][18],A1[26][19],A1[26][20],A1[26][21],A1[26][22],A1[26][23],A1[26][24],A1[26][25],A1[26][26],A1[26][27],A1[27][0],A1[27][1],A1[27][2],A1[27][3],A1[27][4],A1[27][5],A1[27][6],A1[27][7],A1[27][8],A1[27][9],A1[27][10],A1[27][11],A1[27][12],A1[27][13],A1[27][14],A1[27][15],A1[27][16],A1[27][17],A1[27][18],A1[27][19],A1[27][20],A1[27][21],A1[27][22],A1[27][23],A1[27][24],A1[27][25],A1[27][26],A1[27][27]} = A;


        {B1[0][0],B1[0][1],B1[0][2],B1[1][0],B1[1][1],B1[1][2],B1[2][0],B1[2][1],B1[2][2]} = B;

        //initialize to zeros
        
        i = 0;
        j = 0;
        k = 0;

        //initialize to zeros.
        {Res1[0][0],Res1[0][1],Res1[0][2],Res1[0][3],Res1[0][4],Res1[0][5],Res1[0][6],Res1[0][7],Res1[0][8],Res1[0][9],Res1[0][10],Res1[0][11],Res1[0][12],Res1[0][13],Res1[0][14],Res1[0][15],Res1[0][16],Res1[0][17],Res1[0][18],Res1[0][19],Res1[0][20],Res1[0][21],Res1[0][22],Res1[0][23],Res1[0][24],Res1[0][25],Res1[1][0],Res1[1][1],Res1[1][2],Res1[1][3],Res1[1][4],Res1[1][5],Res1[1][6],Res1[1][7],Res1[1][8],Res1[1][9],Res1[1][10],Res1[1][11],Res1[1][12],Res1[1][13],Res1[1][14],Res1[1][15],Res1[1][16],Res1[1][17],Res1[1][18],Res1[1][19],Res1[1][20],Res1[1][21],Res1[1][22],Res1[1][23],Res1[1][24],Res1[1][25],Res1[2][0],Res1[2][1],Res1[2][2],Res1[2][3],Res1[2][4],Res1[2][5],Res1[2][6],Res1[2][7],Res1[2][8],Res1[2][9],Res1[2][10],Res1[2][11],Res1[2][12],Res1[2][13],Res1[2][14],Res1[2][15],Res1[2][16],Res1[2][17],Res1[2][18],Res1[2][19],Res1[2][20],Res1[2][21],Res1[2][22],Res1[2][23],Res1[2][24],Res1[2][25],Res1[3][0],Res1[3][1],Res1[3][2],Res1[3][3],Res1[3][4],Res1[3][5],Res1[3][6],Res1[3][7],Res1[3][8],Res1[3][9],Res1[3][10],Res1[3][11],Res1[3][12],Res1[3][13],Res1[3][14],Res1[3][15],Res1[3][16],Res1[3][17],Res1[3][18],Res1[3][19],Res1[3][20],Res1[3][21],Res1[3][22],Res1[3][23],Res1[3][24],Res1[3][25],Res1[4][0],Res1[4][1],Res1[4][2],Res1[4][3],Res1[4][4],Res1[4][5],Res1[4][6],Res1[4][7],Res1[4][8],Res1[4][9],Res1[4][10],Res1[4][11],Res1[4][12],Res1[4][13],Res1[4][14],Res1[4][15],Res1[4][16],Res1[4][17],Res1[4][18],Res1[4][19],Res1[4][20],Res1[4][21],Res1[4][22],Res1[4][23],Res1[4][24],Res1[4][25],Res1[5][0],Res1[5][1],Res1[5][2],Res1[5][3],Res1[5][4],Res1[5][5],Res1[5][6],Res1[5][7],Res1[5][8],Res1[5][9],Res1[5][10],Res1[5][11],Res1[5][12],Res1[5][13],Res1[5][14],Res1[5][15],Res1[5][16],Res1[5][17],Res1[5][18],Res1[5][19],Res1[5][20],Res1[5][21],Res1[5][22],Res1[5][23],Res1[5][24],Res1[5][25],Res1[6][0],Res1[6][1],Res1[6][2],Res1[6][3],Res1[6][4],Res1[6][5],Res1[6][6],Res1[6][7],Res1[6][8],Res1[6][9],Res1[6][10],Res1[6][11],Res1[6][12],Res1[6][13],Res1[6][14],Res1[6][15],Res1[6][16],Res1[6][17],Res1[6][18],Res1[6][19],Res1[6][20],Res1[6][21],Res1[6][22],Res1[6][23],Res1[6][24],Res1[6][25],Res1[7][0],Res1[7][1],Res1[7][2],Res1[7][3],Res1[7][4],Res1[7][5],Res1[7][6],Res1[7][7],Res1[7][8],Res1[7][9],Res1[7][10],Res1[7][11],Res1[7][12],Res1[7][13],Res1[7][14],Res1[7][15],Res1[7][16],Res1[7][17],Res1[7][18],Res1[7][19],Res1[7][20],Res1[7][21],Res1[7][22],Res1[7][23],Res1[7][24],Res1[7][25],Res1[8][0],Res1[8][1],Res1[8][2],Res1[8][3],Res1[8][4],Res1[8][5],Res1[8][6],Res1[8][7],Res1[8][8],Res1[8][9],Res1[8][10],Res1[8][11],Res1[8][12],Res1[8][13],Res1[8][14],Res1[8][15],Res1[8][16],Res1[8][17],Res1[8][18],Res1[8][19],Res1[8][20],Res1[8][21],Res1[8][22],Res1[8][23],Res1[8][24],Res1[8][25],Res1[9][0],Res1[9][1],Res1[9][2],Res1[9][3],Res1[9][4],Res1[9][5],Res1[9][6],Res1[9][7],Res1[9][8],Res1[9][9],Res1[9][10],Res1[9][11],Res1[9][12],Res1[9][13],Res1[9][14],Res1[9][15],Res1[9][16],Res1[9][17],Res1[9][18],Res1[9][19],Res1[9][20],Res1[9][21],Res1[9][22],Res1[9][23],Res1[9][24],Res1[9][25],Res1[10][0],Res1[10][1],Res1[10][2],Res1[10][3],Res1[10][4],Res1[10][5],Res1[10][6],Res1[10][7],Res1[10][8],Res1[10][9],Res1[10][10],Res1[10][11],Res1[10][12],Res1[10][13],Res1[10][14],Res1[10][15],Res1[10][16],Res1[10][17],Res1[10][18],Res1[10][19],Res1[10][20],Res1[10][21],Res1[10][22],Res1[10][23],Res1[10][24],Res1[10][25],Res1[11][0],Res1[11][1],Res1[11][2],Res1[11][3],Res1[11][4],Res1[11][5],Res1[11][6],Res1[11][7],Res1[11][8],Res1[11][9],Res1[11][10],Res1[11][11],Res1[11][12],Res1[11][13],Res1[11][14],Res1[11][15],Res1[11][16],Res1[11][17],Res1[11][18],Res1[11][19],Res1[11][20],Res1[11][21],Res1[11][22],Res1[11][23],Res1[11][24],Res1[11][25],Res1[12][0],Res1[12][1],Res1[12][2],Res1[12][3],Res1[12][4],Res1[12][5],Res1[12][6],Res1[12][7],Res1[12][8],Res1[12][9],Res1[12][10],Res1[12][11],Res1[12][12],Res1[12][13],Res1[12][14],Res1[12][15],Res1[12][16],Res1[12][17],Res1[12][18],Res1[12][19],Res1[12][20],Res1[12][21],Res1[12][22],Res1[12][23],Res1[12][24],Res1[12][25],Res1[13][0],Res1[13][1],Res1[13][2],Res1[13][3],Res1[13][4],Res1[13][5],Res1[13][6],Res1[13][7],Res1[13][8],Res1[13][9],Res1[13][10],Res1[13][11],Res1[13][12],Res1[13][13],Res1[13][14],Res1[13][15],Res1[13][16],Res1[13][17],Res1[13][18],Res1[13][19],Res1[13][20],Res1[13][21],Res1[13][22],Res1[13][23],Res1[13][24],Res1[13][25],Res1[14][0],Res1[14][1],Res1[14][2],Res1[14][3],Res1[14][4],Res1[14][5],Res1[14][6],Res1[14][7],Res1[14][8],Res1[14][9],Res1[14][10],Res1[14][11],Res1[14][12],Res1[14][13],Res1[14][14],Res1[14][15],Res1[14][16],Res1[14][17],Res1[14][18],Res1[14][19],Res1[14][20],Res1[14][21],Res1[14][22],Res1[14][23],Res1[14][24],Res1[14][25],Res1[15][0],Res1[15][1],Res1[15][2],Res1[15][3],Res1[15][4],Res1[15][5],Res1[15][6],Res1[15][7],Res1[15][8],Res1[15][9],Res1[15][10],Res1[15][11],Res1[15][12],Res1[15][13],Res1[15][14],Res1[15][15],Res1[15][16],Res1[15][17],Res1[15][18],Res1[15][19],Res1[15][20],Res1[15][21],Res1[15][22],Res1[15][23],Res1[15][24],Res1[15][25],Res1[16][0],Res1[16][1],Res1[16][2],Res1[16][3],Res1[16][4],Res1[16][5],Res1[16][6],Res1[16][7],Res1[16][8],Res1[16][9],Res1[16][10],Res1[16][11],Res1[16][12],Res1[16][13],Res1[16][14],Res1[16][15],Res1[16][16],Res1[16][17],Res1[16][18],Res1[16][19],Res1[16][20],Res1[16][21],Res1[16][22],Res1[16][23],Res1[16][24],Res1[16][25],Res1[17][0],Res1[17][1],Res1[17][2],Res1[17][3],Res1[17][4],Res1[17][5],Res1[17][6],Res1[17][7],Res1[17][8],Res1[17][9],Res1[17][10],Res1[17][11],Res1[17][12],Res1[17][13],Res1[17][14],Res1[17][15],Res1[17][16],Res1[17][17],Res1[17][18],Res1[17][19],Res1[17][20],Res1[17][21],Res1[17][22],Res1[17][23],Res1[17][24],Res1[17][25],Res1[18][0],Res1[18][1],Res1[18][2],Res1[18][3],Res1[18][4],Res1[18][5],Res1[18][6],Res1[18][7],Res1[18][8],Res1[18][9],Res1[18][10],Res1[18][11],Res1[18][12],Res1[18][13],Res1[18][14],Res1[18][15],Res1[18][16],Res1[18][17],Res1[18][18],Res1[18][19],Res1[18][20],Res1[18][21],Res1[18][22],Res1[18][23],Res1[18][24],Res1[18][25],Res1[19][0],Res1[19][1],Res1[19][2],Res1[19][3],Res1[19][4],Res1[19][5],Res1[19][6],Res1[19][7],Res1[19][8],Res1[19][9],Res1[19][10],Res1[19][11],Res1[19][12],Res1[19][13],Res1[19][14],Res1[19][15],Res1[19][16],Res1[19][17],Res1[19][18],Res1[19][19],Res1[19][20],Res1[19][21],Res1[19][22],Res1[19][23],Res1[19][24],Res1[19][25],Res1[20][0],Res1[20][1],Res1[20][2],Res1[20][3],Res1[20][4],Res1[20][5],Res1[20][6],Res1[20][7],Res1[20][8],Res1[20][9],Res1[20][10],Res1[20][11],Res1[20][12],Res1[20][13],Res1[20][14],Res1[20][15],Res1[20][16],Res1[20][17],Res1[20][18],Res1[20][19],Res1[20][20],Res1[20][21],Res1[20][22],Res1[20][23],Res1[20][24],Res1[20][25],Res1[21][0],Res1[21][1],Res1[21][2],Res1[21][3],Res1[21][4],Res1[21][5],Res1[21][6],Res1[21][7],Res1[21][8],Res1[21][9],Res1[21][10],Res1[21][11],Res1[21][12],Res1[21][13],Res1[21][14],Res1[21][15],Res1[21][16],Res1[21][17],Res1[21][18],Res1[21][19],Res1[21][20],Res1[21][21],Res1[21][22],Res1[21][23],Res1[21][24],Res1[21][25],Res1[22][0],Res1[22][1],Res1[22][2],Res1[22][3],Res1[22][4],Res1[22][5],Res1[22][6],Res1[22][7],Res1[22][8],Res1[22][9],Res1[22][10],Res1[22][11],Res1[22][12],Res1[22][13],Res1[22][14],Res1[22][15],Res1[22][16],Res1[22][17],Res1[22][18],Res1[22][19],Res1[22][20],Res1[22][21],Res1[22][22],Res1[22][23],Res1[22][24],Res1[22][25],Res1[23][0],Res1[23][1],Res1[23][2],Res1[23][3],Res1[23][4],Res1[23][5],Res1[23][6],Res1[23][7],Res1[23][8],Res1[23][9],Res1[23][10],Res1[23][11],Res1[23][12],Res1[23][13],Res1[23][14],Res1[23][15],Res1[23][16],Res1[23][17],Res1[23][18],Res1[23][19],Res1[23][20],Res1[23][21],Res1[23][22],Res1[23][23],Res1[23][24],Res1[23][25],Res1[24][0],Res1[24][1],Res1[24][2],Res1[24][3],Res1[24][4],Res1[24][5],Res1[24][6],Res1[24][7],Res1[24][8],Res1[24][9],Res1[24][10],Res1[24][11],Res1[24][12],Res1[24][13],Res1[24][14],Res1[24][15],Res1[24][16],Res1[24][17],Res1[24][18],Res1[24][19],Res1[24][20],Res1[24][21],Res1[24][22],Res1[24][23],Res1[24][24],Res1[24][25],Res1[25][0],Res1[25][1],Res1[25][2],Res1[25][3],Res1[25][4],Res1[25][5],Res1[25][6],Res1[25][7],Res1[25][8],Res1[25][9],Res1[25][10],Res1[25][11],Res1[25][12],Res1[25][13],Res1[25][14],Res1[25][15],Res1[25][16],Res1[25][17],Res1[25][18],Res1[25][19],Res1[25][20],Res1[25][21],Res1[25][22],Res1[25][23],Res1[25][24],Res1[25][25]} = 72'd0; 
        

        //Convolution
        for(i=0;i < 26;i=i+1) begin
            for(j=0;j < 26;j=j+1) begin
                Res1[i][j] = Res1[i][j] + A1[i][j] * B1[0][0] + A1[i+1][j] * B1[1][0] + A1[i+2][j] * B1[2][0] + A1[i][j+1] * B1[0][1] + A1[i+1][j+1] * B1[1][1] + A1[i+2][j+1] * B1[2][1] + A1[i][j+2] * B1[0][2] + A1[i+1][j+2] * B1[1][2] + A1[i+2][j+2] * B1[2][2];
            end
        end

        //final output assignment - 3D array to 1D array conversion.            
        Res = {Res1[0][0],Res1[0][1],Res1[0][2],Res1[0][3],Res1[0][4],Res1[0][5],Res1[0][6],Res1[0][7],Res1[0][8],Res1[0][9],Res1[0][10],Res1[0][11],Res1[0][12],Res1[0][13],Res1[0][14],Res1[0][15],Res1[0][16],Res1[0][17],Res1[0][18],Res1[0][19],Res1[0][20],Res1[0][21],Res1[0][22],Res1[0][23],Res1[0][24],Res1[0][25],Res1[1][0],Res1[1][1],Res1[1][2],Res1[1][3],Res1[1][4],Res1[1][5],Res1[1][6],Res1[1][7],Res1[1][8],Res1[1][9],Res1[1][10],Res1[1][11],Res1[1][12],Res1[1][13],Res1[1][14],Res1[1][15],Res1[1][16],Res1[1][17],Res1[1][18],Res1[1][19],Res1[1][20],Res1[1][21],Res1[1][22],Res1[1][23],Res1[1][24],Res1[1][25],Res1[2][0],Res1[2][1],Res1[2][2],Res1[2][3],Res1[2][4],Res1[2][5],Res1[2][6],Res1[2][7],Res1[2][8],Res1[2][9],Res1[2][10],Res1[2][11],Res1[2][12],Res1[2][13],Res1[2][14],Res1[2][15],Res1[2][16],Res1[2][17],Res1[2][18],Res1[2][19],Res1[2][20],Res1[2][21],Res1[2][22],Res1[2][23],Res1[2][24],Res1[2][25],Res1[3][0],Res1[3][1],Res1[3][2],Res1[3][3],Res1[3][4],Res1[3][5],Res1[3][6],Res1[3][7],Res1[3][8],Res1[3][9],Res1[3][10],Res1[3][11],Res1[3][12],Res1[3][13],Res1[3][14],Res1[3][15],Res1[3][16],Res1[3][17],Res1[3][18],Res1[3][19],Res1[3][20],Res1[3][21],Res1[3][22],Res1[3][23],Res1[3][24],Res1[3][25],Res1[4][0],Res1[4][1],Res1[4][2],Res1[4][3],Res1[4][4],Res1[4][5],Res1[4][6],Res1[4][7],Res1[4][8],Res1[4][9],Res1[4][10],Res1[4][11],Res1[4][12],Res1[4][13],Res1[4][14],Res1[4][15],Res1[4][16],Res1[4][17],Res1[4][18],Res1[4][19],Res1[4][20],Res1[4][21],Res1[4][22],Res1[4][23],Res1[4][24],Res1[4][25],Res1[5][0],Res1[5][1],Res1[5][2],Res1[5][3],Res1[5][4],Res1[5][5],Res1[5][6],Res1[5][7],Res1[5][8],Res1[5][9],Res1[5][10],Res1[5][11],Res1[5][12],Res1[5][13],Res1[5][14],Res1[5][15],Res1[5][16],Res1[5][17],Res1[5][18],Res1[5][19],Res1[5][20],Res1[5][21],Res1[5][22],Res1[5][23],Res1[5][24],Res1[5][25],Res1[6][0],Res1[6][1],Res1[6][2],Res1[6][3],Res1[6][4],Res1[6][5],Res1[6][6],Res1[6][7],Res1[6][8],Res1[6][9],Res1[6][10],Res1[6][11],Res1[6][12],Res1[6][13],Res1[6][14],Res1[6][15],Res1[6][16],Res1[6][17],Res1[6][18],Res1[6][19],Res1[6][20],Res1[6][21],Res1[6][22],Res1[6][23],Res1[6][24],Res1[6][25],Res1[7][0],Res1[7][1],Res1[7][2],Res1[7][3],Res1[7][4],Res1[7][5],Res1[7][6],Res1[7][7],Res1[7][8],Res1[7][9],Res1[7][10],Res1[7][11],Res1[7][12],Res1[7][13],Res1[7][14],Res1[7][15],Res1[7][16],Res1[7][17],Res1[7][18],Res1[7][19],Res1[7][20],Res1[7][21],Res1[7][22],Res1[7][23],Res1[7][24],Res1[7][25],Res1[8][0],Res1[8][1],Res1[8][2],Res1[8][3],Res1[8][4],Res1[8][5],Res1[8][6],Res1[8][7],Res1[8][8],Res1[8][9],Res1[8][10],Res1[8][11],Res1[8][12],Res1[8][13],Res1[8][14],Res1[8][15],Res1[8][16],Res1[8][17],Res1[8][18],Res1[8][19],Res1[8][20],Res1[8][21],Res1[8][22],Res1[8][23],Res1[8][24],Res1[8][25],Res1[9][0],Res1[9][1],Res1[9][2],Res1[9][3],Res1[9][4],Res1[9][5],Res1[9][6],Res1[9][7],Res1[9][8],Res1[9][9],Res1[9][10],Res1[9][11],Res1[9][12],Res1[9][13],Res1[9][14],Res1[9][15],Res1[9][16],Res1[9][17],Res1[9][18],Res1[9][19],Res1[9][20],Res1[9][21],Res1[9][22],Res1[9][23],Res1[9][24],Res1[9][25],Res1[10][0],Res1[10][1],Res1[10][2],Res1[10][3],Res1[10][4],Res1[10][5],Res1[10][6],Res1[10][7],Res1[10][8],Res1[10][9],Res1[10][10],Res1[10][11],Res1[10][12],Res1[10][13],Res1[10][14],Res1[10][15],Res1[10][16],Res1[10][17],Res1[10][18],Res1[10][19],Res1[10][20],Res1[10][21],Res1[10][22],Res1[10][23],Res1[10][24],Res1[10][25],Res1[11][0],Res1[11][1],Res1[11][2],Res1[11][3],Res1[11][4],Res1[11][5],Res1[11][6],Res1[11][7],Res1[11][8],Res1[11][9],Res1[11][10],Res1[11][11],Res1[11][12],Res1[11][13],Res1[11][14],Res1[11][15],Res1[11][16],Res1[11][17],Res1[11][18],Res1[11][19],Res1[11][20],Res1[11][21],Res1[11][22],Res1[11][23],Res1[11][24],Res1[11][25],Res1[12][0],Res1[12][1],Res1[12][2],Res1[12][3],Res1[12][4],Res1[12][5],Res1[12][6],Res1[12][7],Res1[12][8],Res1[12][9],Res1[12][10],Res1[12][11],Res1[12][12],Res1[12][13],Res1[12][14],Res1[12][15],Res1[12][16],Res1[12][17],Res1[12][18],Res1[12][19],Res1[12][20],Res1[12][21],Res1[12][22],Res1[12][23],Res1[12][24],Res1[12][25],Res1[13][0],Res1[13][1],Res1[13][2],Res1[13][3],Res1[13][4],Res1[13][5],Res1[13][6],Res1[13][7],Res1[13][8],Res1[13][9],Res1[13][10],Res1[13][11],Res1[13][12],Res1[13][13],Res1[13][14],Res1[13][15],Res1[13][16],Res1[13][17],Res1[13][18],Res1[13][19],Res1[13][20],Res1[13][21],Res1[13][22],Res1[13][23],Res1[13][24],Res1[13][25],Res1[14][0],Res1[14][1],Res1[14][2],Res1[14][3],Res1[14][4],Res1[14][5],Res1[14][6],Res1[14][7],Res1[14][8],Res1[14][9],Res1[14][10],Res1[14][11],Res1[14][12],Res1[14][13],Res1[14][14],Res1[14][15],Res1[14][16],Res1[14][17],Res1[14][18],Res1[14][19],Res1[14][20],Res1[14][21],Res1[14][22],Res1[14][23],Res1[14][24],Res1[14][25],Res1[15][0],Res1[15][1],Res1[15][2],Res1[15][3],Res1[15][4],Res1[15][5],Res1[15][6],Res1[15][7],Res1[15][8],Res1[15][9],Res1[15][10],Res1[15][11],Res1[15][12],Res1[15][13],Res1[15][14],Res1[15][15],Res1[15][16],Res1[15][17],Res1[15][18],Res1[15][19],Res1[15][20],Res1[15][21],Res1[15][22],Res1[15][23],Res1[15][24],Res1[15][25],Res1[16][0],Res1[16][1],Res1[16][2],Res1[16][3],Res1[16][4],Res1[16][5],Res1[16][6],Res1[16][7],Res1[16][8],Res1[16][9],Res1[16][10],Res1[16][11],Res1[16][12],Res1[16][13],Res1[16][14],Res1[16][15],Res1[16][16],Res1[16][17],Res1[16][18],Res1[16][19],Res1[16][20],Res1[16][21],Res1[16][22],Res1[16][23],Res1[16][24],Res1[16][25],Res1[17][0],Res1[17][1],Res1[17][2],Res1[17][3],Res1[17][4],Res1[17][5],Res1[17][6],Res1[17][7],Res1[17][8],Res1[17][9],Res1[17][10],Res1[17][11],Res1[17][12],Res1[17][13],Res1[17][14],Res1[17][15],Res1[17][16],Res1[17][17],Res1[17][18],Res1[17][19],Res1[17][20],Res1[17][21],Res1[17][22],Res1[17][23],Res1[17][24],Res1[17][25],Res1[18][0],Res1[18][1],Res1[18][2],Res1[18][3],Res1[18][4],Res1[18][5],Res1[18][6],Res1[18][7],Res1[18][8],Res1[18][9],Res1[18][10],Res1[18][11],Res1[18][12],Res1[18][13],Res1[18][14],Res1[18][15],Res1[18][16],Res1[18][17],Res1[18][18],Res1[18][19],Res1[18][20],Res1[18][21],Res1[18][22],Res1[18][23],Res1[18][24],Res1[18][25],Res1[19][0],Res1[19][1],Res1[19][2],Res1[19][3],Res1[19][4],Res1[19][5],Res1[19][6],Res1[19][7],Res1[19][8],Res1[19][9],Res1[19][10],Res1[19][11],Res1[19][12],Res1[19][13],Res1[19][14],Res1[19][15],Res1[19][16],Res1[19][17],Res1[19][18],Res1[19][19],Res1[19][20],Res1[19][21],Res1[19][22],Res1[19][23],Res1[19][24],Res1[19][25],Res1[20][0],Res1[20][1],Res1[20][2],Res1[20][3],Res1[20][4],Res1[20][5],Res1[20][6],Res1[20][7],Res1[20][8],Res1[20][9],Res1[20][10],Res1[20][11],Res1[20][12],Res1[20][13],Res1[20][14],Res1[20][15],Res1[20][16],Res1[20][17],Res1[20][18],Res1[20][19],Res1[20][20],Res1[20][21],Res1[20][22],Res1[20][23],Res1[20][24],Res1[20][25],Res1[21][0],Res1[21][1],Res1[21][2],Res1[21][3],Res1[21][4],Res1[21][5],Res1[21][6],Res1[21][7],Res1[21][8],Res1[21][9],Res1[21][10],Res1[21][11],Res1[21][12],Res1[21][13],Res1[21][14],Res1[21][15],Res1[21][16],Res1[21][17],Res1[21][18],Res1[21][19],Res1[21][20],Res1[21][21],Res1[21][22],Res1[21][23],Res1[21][24],Res1[21][25],Res1[22][0],Res1[22][1],Res1[22][2],Res1[22][3],Res1[22][4],Res1[22][5],Res1[22][6],Res1[22][7],Res1[22][8],Res1[22][9],Res1[22][10],Res1[22][11],Res1[22][12],Res1[22][13],Res1[22][14],Res1[22][15],Res1[22][16],Res1[22][17],Res1[22][18],Res1[22][19],Res1[22][20],Res1[22][21],Res1[22][22],Res1[22][23],Res1[22][24],Res1[22][25],Res1[23][0],Res1[23][1],Res1[23][2],Res1[23][3],Res1[23][4],Res1[23][5],Res1[23][6],Res1[23][7],Res1[23][8],Res1[23][9],Res1[23][10],Res1[23][11],Res1[23][12],Res1[23][13],Res1[23][14],Res1[23][15],Res1[23][16],Res1[23][17],Res1[23][18],Res1[23][19],Res1[23][20],Res1[23][21],Res1[23][22],Res1[23][23],Res1[23][24],Res1[23][25],Res1[24][0],Res1[24][1],Res1[24][2],Res1[24][3],Res1[24][4],Res1[24][5],Res1[24][6],Res1[24][7],Res1[24][8],Res1[24][9],Res1[24][10],Res1[24][11],Res1[24][12],Res1[24][13],Res1[24][14],Res1[24][15],Res1[24][16],Res1[24][17],Res1[24][18],Res1[24][19],Res1[24][20],Res1[24][21],Res1[24][22],Res1[24][23],Res1[24][24],Res1[24][25],Res1[25][0],Res1[25][1],Res1[25][2],Res1[25][3],Res1[25][4],Res1[25][5],Res1[25][6],Res1[25][7],Res1[25][8],Res1[25][9],Res1[25][10],Res1[25][11],Res1[25][12],Res1[25][13],Res1[25][14],Res1[25][15],Res1[25][16],Res1[25][17],Res1[25][18],Res1[25][19],Res1[25][20],Res1[25][21],Res1[25][22],Res1[25][23],Res1[25][24],Res1[25][25]};
    end 

endmodule
