 module tb(input wire clk,
    //output wire enable,
    output reg b0,
    output reg b1,
    output reg b2, 
    output reg b3, 
    output reg b4, 
    output reg b5, 
    output reg b6, 
    output reg b7);

    // Inputs
    // Inputs
    reg [3919:0] A;
    reg [26:0] B;
    // Outputs
    reg [5407:0] Res;
    integer i=0;

    // Instantiate the Unit Under Test (UUT)
    sobel_filter filter (
        .A(A), 
        .B(B), 
        .Res(Res)
    );

    initial begin
        // Apply Inputs
        //enable <= 1'b0;
        B <= {3'd1,3'd4,3'd1,3'd0,3'd0,3'd0,-3'd1,-3'd4,-3'd1};
A <= {5'd0,5'd2,5'd1,5'd0,5'd4,5'd2,5'd0,5'd0,5'd2,5'd0,5'd3,5'd9,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd9,5'd0,5'd0,5'd8,5'd0,5'd1,5'd0,5'd0,5'd0,5'd0,5'd5,5'd6,5'd0,5'd0,5'd1,5'd5,5'd3,5'd7,5'd0,5'd11,5'd0,5'd0,5'd4,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd5,5'd7,5'd3,5'd1,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd4,5'd6,5'd0,5'd2,5'd5,5'd9,5'd0,5'd0,5'd14,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd0,5'd3,5'd4,5'd0,5'd0,5'd1,5'd1,5'd4,5'd17,5'd1,5'd0,5'd16,5'd14,5'd0,5'd0,5'd11,5'd0,5'd0,5'd0,5'd14,5'd0,5'd2,5'd0,5'd4,5'd2,5'd0,5'd0,5'd0,5'd0,5'd10,5'd1,5'd0,5'd0,5'd10,5'd5,5'd0,5'd0,5'd8,5'd26,5'd5,5'd23,5'd1,5'd22,5'd28,5'd25,5'd10,5'd0,5'd7,5'd1,5'd0,5'd5,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd2,5'd5,5'd7,5'd5,5'd0,5'd0,5'd14,5'd27,5'd16,5'd31,5'd18,5'd20,5'd31,5'd31,5'd30,5'd25,5'd14,5'd0,5'd3,5'd0,5'd4,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd5,5'd0,5'd0,5'd0,5'd9,5'd30,5'd23,5'd14,5'd17,5'd0,5'd0,5'd0,5'd10,5'd15,5'd31,5'd21,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd1,5'd0,5'd0,5'd1,5'd5,5'd0,5'd0,5'd4,5'd0,5'd3,5'd0,5'd0,5'd9,5'd0,5'd0,5'd0,5'd13,5'd4,5'd0,5'd0,5'd3,5'd0,5'd1,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd0,5'd12,5'd4,5'd3,5'd12,5'd31,5'd16,5'd0,5'd6,5'd1,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd10,5'd0,5'd0,5'd0,5'd4,5'd7,5'd26,5'd19,5'd0,5'd13,5'd5,5'd0,5'd11,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd21,5'd0,5'd0,5'd2,5'd15,5'd12,5'd4,5'd30,5'd19,5'd0,5'd14,5'd0,5'd2,5'd4,5'd6,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd1,5'd26,5'd5,5'd4,5'd31,5'd22,5'd12,5'd4,5'd0,5'd0,5'd0,5'd4,5'd6,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd9,5'd0,5'd30,5'd16,5'd4,5'd13,5'd31,5'd31,5'd30,5'd4,5'd0,5'd0,5'd4,5'd2,5'd0,5'd1,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd22,5'd0,5'd0,5'd15,5'd0,5'd0,5'd2,5'd31,5'd17,5'd10,5'd16,5'd0,5'd0,5'd19,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd7,5'd1,5'd0,5'd2,5'd3,5'd0,5'd8,5'd15,5'd18,5'd31,5'd16,5'd4,5'd0,5'd2,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd8,5'd1,5'd0,5'd11,5'd0,5'd0,5'd0,5'd2,5'd31,5'd31,5'd18,5'd14,5'd0,5'd1,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd2,5'd6,5'd0,5'd0,5'd3,5'd5,5'd0,5'd0,5'd0,5'd1,5'd1,5'd6,5'd0,5'd24,5'd31,5'd4,5'd1,5'd0,5'd2,5'd0,5'd0,5'd0,5'd0,5'd2,5'd5,5'd0,5'd6,5'd20,5'd0,5'd0,5'd1,5'd0,5'd2,5'd6,5'd0,5'd0,5'd0,5'd2,5'd1,5'd0,5'd15,5'd4,5'd19,5'd26,5'd0,5'd17,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd15,5'd0,5'd11,5'd2,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd8,5'd0,5'd23,5'd26,5'd31,5'd0,5'd3,5'd6,5'd0,5'd0,5'd0,5'd0,5'd19,5'd1,5'd0,5'd0,5'd6,5'd0,5'd0,5'd0,5'd8,5'd0,5'd0,5'd3,5'd10,5'd2,5'd0,5'd8,5'd0,5'd3,5'd5,5'd0,5'd15,5'd10,5'd0,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd6,5'd6,5'd0,5'd31,5'd26,5'd0,5'd0,5'd5,5'd13,5'd1,5'd0,5'd0,5'd2,5'd0,5'd2,5'd31,5'd20,5'd10,5'd0,5'd9,5'd0,5'd3,5'd0,5'd0,5'd0,5'd0,5'd16,5'd6,5'd4,5'd0,5'd7,5'd0,5'd0,5'd12,5'd12,5'd7,5'd0,5'd11,5'd8,5'd0,5'd28,5'd2,5'd26,5'd17,5'd24,5'd13,5'd0,5'd0,5'd10,5'd3,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd0,5'd0,5'd20,5'd8,5'd30,5'd6,5'd31,5'd31,5'd11,5'd26,5'd30,5'd20,5'd7,5'd17,5'd23,5'd5,5'd3,5'd1,5'd4,5'd2,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd3,5'd0,5'd0,5'd4,5'd17,5'd18,5'd30,5'd1,5'd21,5'd7,5'd11,5'd19,5'd30,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0};
    end
    
     
    
    //if(Res) begin    
        always@(posedge clk) begin
            {b7, b6, b5, b4, b3, b2, b1, b0} <= Res[i+7:i];
            i <= i+8;
            //if(i==5400) begin
            //    send_start = 0'b1;
            //end
        end
    //end

endmodule
